`include "pc_control.v"
module pc_control_tb();
    
    
endmodule